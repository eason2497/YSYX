module ps2_keyboard(
	input clk,
	input resetn,
	input ps2_clk,
	input ps2_data,
	output reg [3:0] press,
	output reg [3:0] bcd1,
	output reg [3:0] bcd2
);

    reg [9:0] buffer;        // ps2_data bits
    reg [3:0] count;  // count ps2_data bits
    reg [2:0] ps2_clk_sync;
    reg pressing;
    initial 
    begin
    press = 4'b0;
    pressing = 0;
    end    
    
    always @(posedge clk) begin
        ps2_clk_sync <=  {ps2_clk_sync[1:0],ps2_clk};
    end

    wire sampling = ps2_clk_sync[2] & ~ps2_clk_sync[1];
    always @(posedge clk) begin
        if (resetn == 0) begin // reset
            count <= 0;
        end
        else begin
            if (sampling) begin
	      press <= press + 4'b1;
	      if (count == 4'd10) begin
                if ((buffer[0] == 0) &&  // start bit
                    (ps2_data)       &&  // stop bit
                    (^buffer[9:1])) begin      // odd  parity
                    $display("receive %x", buffer[8:1]);
		    bcd1 <= buffer[8:5];
		    bcd2 <= buffer[4:1];
                end
                count <= 0;     // for next
              end else begin
                buffer[count] <= ps2_data;  // store ps2_data
                count <= count + 3'b1;
              end
            end
        end
    end

endmodule
